.title KonCEPT LC-resonanskrets

* Detta är en parallell LC-resonanskrets som kan användas
* för att demonstrera resonans vid en specifik frekvens.

* Strömkälla: 1 mA AC
Iin input 0 AC 1m

* Induktor: 100 uH
L1 input 0 100u

* Kondensator: 100 pF
C1 input 0 100p

* Resistor för förluster: 1 kOhm
R1 input 0 1k

* AC-analys från 100 kHz till 10 MHz med 100 punkter per dekad
.ac dec 100 100k 10meg

.save V(input)
.plot ac V(input)
.hardcopy
.end
